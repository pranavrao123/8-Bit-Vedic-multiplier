module Subtractor(
    input [7:0] A, B,
    output [7:0] result
);
    assign result = A - B;
endmodule
